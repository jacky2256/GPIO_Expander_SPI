module spi2apb_bridge(input );



endmodule